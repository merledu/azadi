package brq_pkg;
    


endpackage
