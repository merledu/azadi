package azadi_pkg;
    


endpackage
